module transmitter(
	);
endmodule
