module transmitter(
	
		);
endmodule
