module synchro(
	);
endmodule
