module uart(
	input i_rst,
	input i_clk,
	output[4:0] o_address,
	output o_read,
	input[31:0] i_readdata,
	output o_write,
	output[31:0] o_writedata,
	input i_waitrequest,

	input[7:0] i_char,
	output[15:0] o_char
	);

//parameters

//logics

//combinational

//sequential

endmodule
