module sdram(
	);

endmodule
