module top(
	
		);
endmodule
